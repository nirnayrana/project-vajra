module vajra_caravel_soc (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire net2;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net3;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net4;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net40;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net41;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net42;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net1;

 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_2 (.LO(net2));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_3 (.LO(net3));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_4 (.LO(net4));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_5 (.LO(net5));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_6 (.LO(net6));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_7 (.LO(net7));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_8 (.LO(net8));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_9 (.LO(net9));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_10 (.LO(net10));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_11 (.LO(net11));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_12 (.LO(net12));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_13 (.LO(net13));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_14 (.LO(net14));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_15 (.LO(net15));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_16 (.LO(net16));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_17 (.LO(net17));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_18 (.LO(net18));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_19 (.LO(net19));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_20 (.LO(net20));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_21 (.LO(net21));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_22 (.LO(net22));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_23 (.LO(net23));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_24 (.LO(net24));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_25 (.LO(net25));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_26 (.LO(net26));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_27 (.LO(net27));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_28 (.LO(net28));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_29 (.LO(net29));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_30 (.LO(net30));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_31 (.LO(net31));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_32 (.LO(net32));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_33 (.LO(net33));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_34 (.LO(net34));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_35 (.LO(net35));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_36 (.LO(net36));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_37 (.LO(net37));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_38 (.LO(net38));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_39 (.LO(net39));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_40 (.LO(net40));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_41 (.LO(net41));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_42 (.LO(net42));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_43 (.LO(net43));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_44 (.LO(net44));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_45 (.LO(net45));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_46 (.LO(net46));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_47 (.LO(net47));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_69 (.LO(net69));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_70 (.LO(net70));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_71 (.LO(net71));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_72 (.LO(net72));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_73 (.LO(net73));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_74 (.LO(net74));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_75 (.LO(net75));
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_76 (.LO(net76));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_6 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_572 ();
 sky130_fd_sc_hd__decap_3 PHY_573 ();
 sky130_fd_sc_hd__decap_3 PHY_574 ();
 sky130_fd_sc_hd__decap_3 PHY_575 ();
 sky130_fd_sc_hd__decap_3 PHY_576 ();
 sky130_fd_sc_hd__decap_3 PHY_577 ();
 sky130_fd_sc_hd__decap_3 PHY_578 ();
 sky130_fd_sc_hd__decap_3 PHY_579 ();
 sky130_fd_sc_hd__decap_3 PHY_580 ();
 sky130_fd_sc_hd__decap_3 PHY_581 ();
 sky130_fd_sc_hd__decap_3 PHY_582 ();
 sky130_fd_sc_hd__decap_3 PHY_583 ();
 sky130_fd_sc_hd__decap_3 PHY_584 ();
 sky130_fd_sc_hd__decap_3 PHY_585 ();
 sky130_fd_sc_hd__decap_3 PHY_586 ();
 sky130_fd_sc_hd__decap_3 PHY_587 ();
 sky130_fd_sc_hd__decap_3 PHY_588 ();
 sky130_fd_sc_hd__decap_3 PHY_589 ();
 sky130_fd_sc_hd__decap_3 PHY_590 ();
 sky130_fd_sc_hd__decap_3 PHY_591 ();
 sky130_fd_sc_hd__decap_3 PHY_592 ();
 sky130_fd_sc_hd__decap_3 PHY_593 ();
 sky130_fd_sc_hd__decap_3 PHY_594 ();
 sky130_fd_sc_hd__decap_3 PHY_595 ();
 sky130_fd_sc_hd__decap_3 PHY_596 ();
 sky130_fd_sc_hd__decap_3 PHY_597 ();
 sky130_fd_sc_hd__decap_3 PHY_598 ();
 sky130_fd_sc_hd__decap_3 PHY_599 ();
 sky130_fd_sc_hd__decap_3 PHY_600 ();
 sky130_fd_sc_hd__decap_3 PHY_601 ();
 sky130_fd_sc_hd__decap_3 PHY_602 ();
 sky130_fd_sc_hd__decap_3 PHY_603 ();
 sky130_fd_sc_hd__decap_3 PHY_604 ();
 sky130_fd_sc_hd__decap_3 PHY_605 ();
 sky130_fd_sc_hd__decap_3 PHY_606 ();
 sky130_fd_sc_hd__decap_3 PHY_607 ();
 sky130_fd_sc_hd__decap_3 PHY_608 ();
 sky130_fd_sc_hd__decap_3 PHY_609 ();
 sky130_fd_sc_hd__decap_3 PHY_610 ();
 sky130_fd_sc_hd__decap_3 PHY_611 ();
 sky130_fd_sc_hd__decap_3 PHY_612 ();
 sky130_fd_sc_hd__decap_3 PHY_613 ();
 sky130_fd_sc_hd__decap_3 PHY_614 ();
 sky130_fd_sc_hd__decap_3 PHY_615 ();
 sky130_fd_sc_hd__decap_3 PHY_616 ();
 sky130_fd_sc_hd__decap_3 PHY_617 ();
 sky130_fd_sc_hd__decap_3 PHY_618 ();
 sky130_fd_sc_hd__decap_3 PHY_619 ();
 sky130_fd_sc_hd__decap_3 PHY_620 ();
 sky130_fd_sc_hd__decap_3 PHY_621 ();
 sky130_fd_sc_hd__decap_3 PHY_622 ();
 sky130_fd_sc_hd__decap_3 PHY_623 ();
 sky130_fd_sc_hd__decap_3 PHY_624 ();
 sky130_fd_sc_hd__decap_3 PHY_625 ();
 sky130_fd_sc_hd__decap_3 PHY_626 ();
 sky130_fd_sc_hd__decap_3 PHY_627 ();
 sky130_fd_sc_hd__decap_3 PHY_628 ();
 sky130_fd_sc_hd__decap_3 PHY_629 ();
 sky130_fd_sc_hd__decap_3 PHY_630 ();
 sky130_fd_sc_hd__decap_3 PHY_631 ();
 sky130_fd_sc_hd__decap_3 PHY_632 ();
 sky130_fd_sc_hd__decap_3 PHY_633 ();
 sky130_fd_sc_hd__decap_3 PHY_634 ();
 sky130_fd_sc_hd__decap_3 PHY_635 ();
 sky130_fd_sc_hd__decap_3 PHY_636 ();
 sky130_fd_sc_hd__decap_3 PHY_637 ();
 sky130_fd_sc_hd__decap_3 PHY_638 ();
 sky130_fd_sc_hd__decap_3 PHY_639 ();
 sky130_fd_sc_hd__decap_3 PHY_640 ();
 sky130_fd_sc_hd__decap_3 PHY_641 ();
 sky130_fd_sc_hd__decap_3 PHY_642 ();
 sky130_fd_sc_hd__decap_3 PHY_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_11659 ();
 sky130_fd_sc_hd__conb_1 vajra_caravel_soc_1 (.LO(net1));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_846 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1238 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1250 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1425 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1434 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1485 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_1650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1681 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1700 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1877 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_1889 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_1896 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_131_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_132_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_134_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_136_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_136_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_137_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_138_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_138_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_139_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_140_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_141_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_142_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_143_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_144_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_145_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_147_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_148_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_149_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_149_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_150_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_151_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_153_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_154_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_155_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_157_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_157_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_157_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_158_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_158_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_158_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_159_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_159_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_159_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_160_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_160_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_160_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_160_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_160_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_160_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_161_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_161_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_161_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_162_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_162_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_162_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_162_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_163_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_163_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_163_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_164_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_164_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_164_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_165_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_165_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_165_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_166_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_166_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_166_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_166_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_167_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_167_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_168_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_168_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_168_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_168_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_169_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_170_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_170_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_170_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_170_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_171_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_171_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_171_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_171_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_172_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_172_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_172_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_172_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_173_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_173_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_173_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_174_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_174_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_174_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_174_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_175_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_175_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_175_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_176_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_176_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_176_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_176_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_177_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_177_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_177_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_178_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_178_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_178_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_178_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_179_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_179_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_179_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_180_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_180_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_180_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_180_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_181_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_181_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_182_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_182_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_182_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_182_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_183_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_183_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_184_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_184_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_184_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_184_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_185_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_185_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_186_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_186_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_186_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_187_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_187_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_187_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_188_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_188_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_188_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_188_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_189_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_189_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_190_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_190_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_190_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_190_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_191_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_191_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_192_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_192_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_192_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_193_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_193_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_193_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_194_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_194_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_194_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_194_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_195_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_195_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_196_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_196_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_196_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_196_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_197_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_197_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_197_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_198_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_198_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_198_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_198_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_199_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_199_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_199_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_200_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_200_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_200_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_200_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_201_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_201_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_201_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_202_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_202_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_202_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_202_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_203_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_203_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_203_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_204_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_204_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_204_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_205_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_205_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_205_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_206_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_206_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_206_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_206_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_207_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_207_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_208_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_208_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_208_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_208_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_209_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_209_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_210_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_210_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_211_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_211_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_211_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_212_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_212_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_212_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_212_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_213_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_213_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_213_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_214_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_214_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_214_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_215_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_215_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_215_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_216_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_216_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_216_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_216_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_217_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_217_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_218_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_218_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_218_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_218_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_219_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_219_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_219_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_219_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_220_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_220_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_220_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_220_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_221_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_221_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_221_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_221_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_222_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_222_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_222_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_222_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_223_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_223_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_224_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_224_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_224_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_224_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_225_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_226_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_226_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_226_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_226_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_227_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_227_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_227_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_228_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_228_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_228_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_228_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_229_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_229_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_230_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_230_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_230_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_230_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_231_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_231_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_232_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_232_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_232_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_233_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_233_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_233_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_234_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_234_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_234_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_234_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_235_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_235_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_235_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_236_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_236_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_236_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_236_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_237_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_237_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_238_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_238_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_238_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_239_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_239_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_239_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_240_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_240_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_240_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_240_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_241_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_241_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_242_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_242_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_242_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_242_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_242_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_242_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_243_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_243_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_243_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_244_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_244_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_244_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_245_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_245_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_245_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_245_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_246_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_246_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_246_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_246_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_247_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_247_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_248_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_248_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_248_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_249_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_249_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_249_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_250_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_250_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_250_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_250_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_251_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_251_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_251_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_252_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_252_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_252_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_252_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_253_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_254_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_254_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_254_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_254_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_255_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_255_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_255_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_256_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_256_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_256_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_257_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_257_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_257_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_258_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_258_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_258_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_258_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_259_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_259_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_260_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_260_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_260_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_260_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_261_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_261_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_262_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_262_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_262_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_262_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_263_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_263_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_264_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_264_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_264_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_264_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_265_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_265_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_266_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_266_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_266_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_266_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_266_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_266_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_267_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_267_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_267_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_268_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_268_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_268_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_268_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_269_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_269_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_269_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_269_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_270_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_270_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_270_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_270_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_271_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_271_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_271_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_272_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_272_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_272_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_272_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_273_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_273_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_274_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_274_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_274_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_274_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_275_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_275_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_275_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_276_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_276_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_276_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_276_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_277_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_277_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_277_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_277_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_278_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_278_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_278_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_278_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_279_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_279_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_280_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_280_1913 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_280_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_281_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_282_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_282_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_282_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_282_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_283_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_283_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_283_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_284_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_284_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_284_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_284_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_285_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_285_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_285_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_286_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_286_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_286_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_286_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_287_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_287_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_287_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_287_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_288_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_288_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_288_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_288_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_289_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_289_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_289_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_289_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_290_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_290_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_290_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_290_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_291_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_291_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_292_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_292_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_292_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_292_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_293_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_293_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_293_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_294_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_294_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_294_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_294_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_295_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_295_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_295_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_295_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_296_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_296_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_296_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_296_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_297_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_297_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_297_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_298_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_298_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_298_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_298_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_299_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_299_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_299_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_300_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_300_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_300_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_300_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_301_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_301_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_301_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_301_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_302_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_302_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_302_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_302_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_303_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_303_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_304_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_304_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_304_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_304_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_305_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_305_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_305_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_305_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_306_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_306_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_306_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_306_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_307_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_307_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_307_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_308_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_308_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_308_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_308_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_309_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_310_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_310_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_310_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_310_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_311_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_311_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_311_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_311_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_312_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_312_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_312_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_312_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_313_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_313_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_313_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_314_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_314_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_314_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_314_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_315_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_315_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_315_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_316_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_316_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_316_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_316_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_317_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_317_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_317_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_317_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_318_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_318_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_318_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_318_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1493 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_319_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_319_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_320_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_320_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_320_1913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_320_1925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_321_1217 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_1510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1537 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1793 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_321_1873 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1882 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1894 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_321_1902 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321_1905 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_321_1917 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_321_1925 ();
 assign io_oeb[0] = net1;
 assign io_oeb[10] = net11;
 assign io_oeb[11] = net12;
 assign io_oeb[12] = net13;
 assign io_oeb[13] = net14;
 assign io_oeb[14] = net15;
 assign io_oeb[15] = net16;
 assign io_oeb[16] = net17;
 assign io_oeb[17] = net18;
 assign io_oeb[18] = net19;
 assign io_oeb[19] = net20;
 assign io_oeb[1] = net2;
 assign io_oeb[20] = net21;
 assign io_oeb[21] = net22;
 assign io_oeb[22] = net23;
 assign io_oeb[23] = net24;
 assign io_oeb[24] = net25;
 assign io_oeb[25] = net26;
 assign io_oeb[26] = net27;
 assign io_oeb[27] = net28;
 assign io_oeb[28] = net29;
 assign io_oeb[29] = net30;
 assign io_oeb[2] = net3;
 assign io_oeb[30] = net31;
 assign io_oeb[31] = net32;
 assign io_oeb[32] = net33;
 assign io_oeb[33] = net34;
 assign io_oeb[34] = net35;
 assign io_oeb[35] = net36;
 assign io_oeb[36] = net37;
 assign io_oeb[37] = net38;
 assign io_oeb[3] = net4;
 assign io_oeb[4] = net5;
 assign io_oeb[5] = net6;
 assign io_oeb[6] = net7;
 assign io_oeb[7] = net8;
 assign io_oeb[8] = net9;
 assign io_oeb[9] = net10;
 assign io_out[0] = net39;
 assign io_out[10] = net49;
 assign io_out[11] = net50;
 assign io_out[12] = net51;
 assign io_out[13] = net52;
 assign io_out[14] = net53;
 assign io_out[15] = net54;
 assign io_out[16] = net55;
 assign io_out[17] = net56;
 assign io_out[18] = net57;
 assign io_out[19] = net58;
 assign io_out[1] = net40;
 assign io_out[20] = net59;
 assign io_out[21] = net60;
 assign io_out[22] = net61;
 assign io_out[23] = net62;
 assign io_out[24] = net63;
 assign io_out[25] = net64;
 assign io_out[26] = net65;
 assign io_out[27] = net66;
 assign io_out[28] = net67;
 assign io_out[29] = net68;
 assign io_out[2] = net41;
 assign io_out[30] = net69;
 assign io_out[31] = net70;
 assign io_out[32] = net71;
 assign io_out[33] = net72;
 assign io_out[34] = net73;
 assign io_out[35] = net74;
 assign io_out[36] = net75;
 assign io_out[37] = net76;
 assign io_out[3] = net42;
 assign io_out[4] = net43;
 assign io_out[5] = net44;
 assign io_out[6] = net45;
 assign io_out[7] = net46;
 assign io_out[8] = net47;
 assign io_out[9] = net48;
endmodule
